// -----------------------------------------------------------------------------
// 模块名称：adc_capture
// 功能描述：
//    采集AD9248复用模式下的双通道数据（A/B通道共用一组数据线），
//    在时钟上升沿采集A通道数据，在时钟下降沿采集B通道数据，
//    并完成无符号转有符号补码转换。
//    输出带符号（signed）的采样数据，便于后续与IP核（如FFT、FIR）对接。
// 端口说明：
//    clk：              时钟
//    data：             14位复用数据输入（A/B通道）
//    a_data_signed：    A通道已转换的有符号输出
//    b_data_signed：    B通道已转换的有符号输出
// -----------------------------------------------------------------------------

module adc_capture (
    input  wire              clk,             // AD采样时钟
    input  wire [13:0]       data_in,            // 14位复用ADC数据输入

    output reg [27:0] data_out
);
    // =========================================================================
    // 采样并编码转换：在各自ADC采样时钟沿完成无符号数 [0,2^14-1] -→ [-2^13,2^13-1]有符号补码
    // =========================================================================

    // 时钟上升沿采样A通道
    always @(posedge clk) begin
        // 采样数据减去2^13，区间平移[0,16383] -→ [-8192,8191]，变为补码形式
        data_out[27:14] <= $signed(data_in) - 14'sd8192;
    end

    // 时钟下降沿采样B通道
    always @(negedge clk) begin
        data_out[13:0] <= $signed(data_in) - 14'sd8192;
    end
endmodule